interface moka_rv32i_sc_if(input clk);
    logic rstn;
    logic en;
endinterface